// 4-bit ones counter circuit
module onescount_4bit(A, O);
  input [3:0] A;
  output [2:0] O;
  reg [2:0] count_ones; 
  integer idx;

  always_comb begin
    count_ones = 0;
    for( idx=0; idx<4; idx=idx+1) begin
      count_ones = count_ones + A[idx];
    end
  end

  assign O = count_ones;

endmodule
